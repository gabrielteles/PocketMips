--Acad�micos:
--Cauan Gama
--Gabriel Teles
--Professor: Ricardo
--Ci�ncia da Computa��o - UFMS 
entity AC is 
end entity;

architecture comportamental of AC is
begin
end architecture;
