entity BC is 
end entity;
architecture comportamental of BC is
end architecture;
