entity AC is 
end entity;

architecture comportamental of AC is
end architecture;
