--Acad�micos:
--Cauan Gama
--Gabriel Teles
--Professor: Ricardo
--Ci�ncia da Computa��o - UFMS 
entity BC is 
end entity;
architecture comportamental of BC is
end architecture;
