entity clock_generator is
	port(
		Halt : in bit;-- parada
		Clk  : out bit;-- clock
		
end entity;
